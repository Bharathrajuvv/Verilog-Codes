// Design code for Not gate 
module notgate (input a,output b);
  not (b,a);
endmodule
